`default_nettype none // prevents system from inferring an undeclared logic (good practice)
 
module top_level(
  input wire sysclk, //crystal reference clock
  input wire [1:0] sw, //all 16 input slide switches
  input wire [3:0] btn, //all four momentary button switches
  output logic [1:0] led, //16 green output LEDs (located right above switches)
//  output logic [2:0] rgb0, //rgb led
 // output logic [2:0] rgb1, //rgb led
  output logic [2:0] hdmi_tx_p, //hdmi output signals (positives) (blue, green, red)
  output logic [2:0] hdmi_tx_n, //hdmi output signals (negatives) (blue, green, red)
  output logic hdmi_clk_p, hdmi_clk_n //differential hdmi clock
  );
 
  assign led = sw; //to verify the switch values
  //shut up those rgb LEDs (active high):
//  assign rgb1= 0;
 // assign rgb0 = 0;
 
  //have btn[0] control system reset
  logic sys_rst;
  assign sys_rst = btn[0]; //reset is btn[0]
  logic game_rst;
  assign game_rst = btn[1]; //reset is btn[1]
 
  logic clk_pixel, clk_5x; //clock lines    
  logic locked; //locked signal (we'll leave unused but still hook it up)
 

      
   clk_wiz_0 clk_inst
  (
  // Clock out ports  
  .clk_out1(clk_pixel),
  .clk_out2(clk_5x),
  // Status and control signals               
  .reset(0), 
  .locked(locked),
 // Clock in ports
  .clk_in1(sysclk)
  );
      
      
      
 
  logic [10:0] hcount; //hcount of system!
  logic [9:0] vcount; //vcount of system!
  logic hor_sync; //horizontal sync signal
  logic vert_sync; //vertical sync signal
  logic active_draw; //ative draw! 1 when in drawing region.0 in blanking/sync
  logic new_frame; //one cycle active indicator of new frame of info!
  logic [5:0] frame_count; //0 to 59 then rollover frame counter
 
 
  video_sig_generator mvg(
      .pixel_clk_in(clk_pixel),
      .rst_in(sys_rst),
      .x(hcount),
      .y(vcount),
      .vs_out(vert_sync),
      .hs_out(hor_sync),
      .ad_out(active_draw),
      .nf_out(new_frame),
     .fc_out(frame_count)
      );
 
  logic [7:0] red, green, blue; //red green and blue pixel values for output
  logic [7:0] tp_r, tp_g, tp_b; //color values as generated by test_pattern module
  logic [7:0] pg_r, pg_g, pg_b;//color values as generated by pong game(part 2)
 
  //comment out in checkoff 1 once you know you have your video pipeline working:
  //these three colors should be a nice pink (6.205 sidebar) color on full screen .

 
  //uncomment the test pattern generator for the latter portion of part 1
  //and use it to drive tp_r,g, and b once you know that your video
  //pipeline is working (by seeing the 6.205 pink color)
  
  test_pattern_generator mtpg(
      .sel_in(sw[1:0]),
      .hcount_in(hcount),
      .vcount_in(vcount),
      .red_out(tp_r),
      .green_out(tp_g),
      .blue_out(tp_b));
  
 
  pong my_pong (
      .pixel_clk_in(clk_pixel),
      .rst_in(game_rst),
      .control_in({clean_b3,clean_b2}),
      .puck_speed_in(4'b0001),
      .paddle_speed_in(4'b0001),
      .nf_in(new_frame),
      .hcount_in(hcount),
      .vcount_in(vcount),
      .red_out(pg_r),
      .green_out(pg_g),
      .blue_out(pg_b));
  
 
  always_comb begin
    if (~sw[1])begin //if switch 3 switched use shapes signal from part 2, else defaults
      red = tp_r;
      green = tp_g;
      blue = tp_b;
    end else begin
      red = pg_r;
      green = pg_g;
      blue = pg_b;
    end
  end
 
  logic [9:0] tmds_10b [0:2]; //output of each TMDS encoder!
  logic tmds_signal [2:0]; //output of each TMDS serializer!
 
  logic clean_b3;//Filtered button 3 value 
  logic clean_b2;//Filtered button 3 value 


 debounce debounce_btn2(
    .clk(clk_pixel),
    .reset(sys_rst),
    .dirty_in(btn(2)),
    .clean_out(clean_b2)
 );
 debounce debounce_btn3(
    .clk(clk_pixel),
    .reset(sys_rst),
    .dirty_in(btn(3)),
    .clean_out(clean_b3)
 );
 
  tmds_encoder tmds_red(
      .clk_in(clk_pixel),
      .rst_in(sys_rst),
      .data_in(red),
      .control_in(2'b0),
      .ve_in(active_draw),
      .tmds_out(tmds_10b[2]));
 
 tmds_encoder tmds_green(
    .clk_in(clk_pixel),
    .rst_in(sys_rst),
    .data_in(green),
    .control_in(2'b0),
    .ve_in(active_draw),
    .tmds_out(tmds_10b[1]));

tmds_encoder tmds_blue(
    .clk_in(clk_pixel),
    .rst_in(sys_rst),
    .data_in(blue),
    .control_in({vert_sync, hor_sync}), // {vsync, hsync}
    .ve_in(active_draw), // only send data during active draw
    .tmds_out(tmds_10b[0]));
 
  //three tmds_serializers (blue, green, red):
  //MISSING: two more serializers for the green and blue tmds signals.
  tmds_serializer red_ser(
      .clk_pixel_in(clk_pixel),
      .clk_5x_in(clk_5x),
      .rst_in(sys_rst),
      .tmds_in(tmds_10b[2]),
      .tmds_out(tmds_signal[2]));
      
      
      tmds_serializer green_ser(
    .clk_pixel_in(clk_pixel),
    .clk_5x_in(clk_5x),
    .rst_in(sys_rst),
    .tmds_in(tmds_10b[1]),
    .tmds_out(tmds_signal[1]));

tmds_serializer blue_ser(
    .clk_pixel_in(clk_pixel),
    .clk_5x_in(clk_5x),
    .rst_in(sys_rst),
    .tmds_in(tmds_10b[0]),
    .tmds_out(tmds_signal[0]));

 
  //output buffers generating differential signals:
  //three for the r,g,b signals and one that is at the pixel clock rate
  //the HDMI receivers use recover logic coupled with the control signals asserted
  //during blanking and sync periods to synchronize their faster bit clocks off
  //of the slower pixel clock (so they can recover a clock of about 742.5 MHz from
  //the slower 74.25 MHz clock)
  OBUFDS OBUFDS_blue (.I(tmds_signal[0]), .O(hdmi_tx_p[0]), .OB(hdmi_tx_n[0]));
  OBUFDS OBUFDS_green(.I(tmds_signal[1]), .O(hdmi_tx_p[1]), .OB(hdmi_tx_n[1]));
  OBUFDS OBUFDS_red  (.I(tmds_signal[2]), .O(hdmi_tx_p[2]), .OB(hdmi_tx_n[2]));
  OBUFDS OBUFDS_clock(.I(clk_pixel), .O(hdmi_clk_p), .OB(hdmi_clk_n));
 
endmodule // top_level
`default_nettype wire